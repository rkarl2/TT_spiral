`default_nettype none
module hypCal (
	input wire [9:0] x_pos,
	input wire [9:0] y_pos,
	input wire clk, rst,
	output reg [3:0] r_sqroot
);
wire [12:0] xy_pos;
wire _unused = &{x_pos[1:0],y_pos[1:0]};

wire  [6:0] norm_x = (x_pos[9] == 1'b0) ? x_pos[8:2] : ~(x_pos[8:2]);
wire  [6:0] norm_y = (y_pos[9] == 1'b0) ? y_pos[8:2] : ~(y_pos[8:2]);

reg [6:0]mutlReg;
reg stateCheck;
wire [12:0]multSignal = mutlReg*mutlReg;
reg[12:0] multX, multY;
always @(posedge clk) begin
	if (rst) begin
		mutlReg <= 7'h00;
		stateCheck <= 'b0;
	end else begin
		if (stateCheck == 'b0) begin
			multY <=multSignal;
			mutlReg <= norm_x;
			stateCheck <= 'b1;
		end else begin
			multX <=multSignal;
			mutlReg <= norm_y;
			stateCheck <= 'b0;
		end
	end
end
		

//assign xy_pos = (norm_y[8:2]*norm_y[8:2] + norm_x[8:2]*norm_x[8:2]) >> 6;
assign xy_pos = (multX + multY) >> 6;
always @(xy_pos) begin
	case(xy_pos)
		'h00 : r_sqroot <= 'h0;
		'h01 : r_sqroot <= 'h3;
		'h02 : r_sqroot <= 'h5;
		'h03 : r_sqroot <= 'h6;
		'h04 : r_sqroot <= 'h7;
		'h05 : r_sqroot <= 'h8;
		'h06 : r_sqroot <= 'h8;
		'h07 : r_sqroot <= 'h9;
		'h08 : r_sqroot <= 'ha;
		'h09 : r_sqroot <= 'ha;
		'h0a : r_sqroot <= 'hb;
		'h0b : r_sqroot <= 'hc;
		'h0c : r_sqroot <= 'hc;
		'h0d : r_sqroot <= 'hd;
		'h0e : r_sqroot <= 'hd;
		'h0f : r_sqroot <= 'he;
		'h10 : r_sqroot <= 'he;
		'h11 : r_sqroot <= 'he;
		'h12 : r_sqroot <= 'hf;
		'h13 : r_sqroot <= 'hf;
		'h14 : r_sqroot <= 'h0;
		'h15 : r_sqroot <= 'h0;
		'h16 : r_sqroot <= 'h0;
		'h17 : r_sqroot <= 'h1;
		'h18 : r_sqroot <= 'h1;
		'h19 : r_sqroot <= 'h2;
		'h1a : r_sqroot <= 'h2;
		'h1b : r_sqroot <= 'h2;
		'h1c : r_sqroot <= 'h3;
		'h1d : r_sqroot <= 'h3;
		'h1e : r_sqroot <= 'h3;
		'h1f : r_sqroot <= 'h4;
		'h20 : r_sqroot <= 'h4;
		'h21 : r_sqroot <= 'h4;
		'h22 : r_sqroot <= 'h5;
		'h23 : r_sqroot <= 'h5;
		'h24 : r_sqroot <= 'h5;
		'h25 : r_sqroot <= 'h6;
		'h26 : r_sqroot <= 'h6;
		'h27 : r_sqroot <= 'h6;
		'h28 : r_sqroot <= 'h6;
		'h29 : r_sqroot <= 'h7;
		'h2a : r_sqroot <= 'h7;
		'h2b : r_sqroot <= 'h7;
		'h2c : r_sqroot <= 'h8;
		'h2d : r_sqroot <= 'h8;
		'h2e : r_sqroot <= 'h8;
		'h2f : r_sqroot <= 'h8;
		'h30 : r_sqroot <= 'h9;
		'h31 : r_sqroot <= 'h9;
		'h32 : r_sqroot <= 'h9;
		'h33 : r_sqroot <= 'h9;
		'h34 : r_sqroot <= 'ha;
		'h35 : r_sqroot <= 'ha;
		'h36 : r_sqroot <= 'ha;
		'h37 : r_sqroot <= 'ha;
		'h38 : r_sqroot <= 'hb;
		'h39 : r_sqroot <= 'hb;
		'h3a : r_sqroot <= 'hb;
		'h3b : r_sqroot <= 'hb;
		'h3c : r_sqroot <= 'hc;
		'h3d : r_sqroot <= 'hc;
		'h3e : r_sqroot <= 'hc;
		'h3f : r_sqroot <= 'hc;
		'h40 : r_sqroot <= 'hc;
		'h41 : r_sqroot <= 'hd;
		'h42 : r_sqroot <= 'hd;
		'h43 : r_sqroot <= 'hd;
		'h44 : r_sqroot <= 'hd;
		'h45 : r_sqroot <= 'he;
		'h46 : r_sqroot <= 'he;
		'h47 : r_sqroot <= 'he;
		'h48 : r_sqroot <= 'he;
		'h49 : r_sqroot <= 'he;
		'h4a : r_sqroot <= 'hf;
		'h4b : r_sqroot <= 'hf;
		'h4c : r_sqroot <= 'hf;
		'h4d : r_sqroot <= 'hf;
		'h4e : r_sqroot <= 'hf;
		'h4f : r_sqroot <= 'h0;
		'h50 : r_sqroot <= 'h0;
		'h51 : r_sqroot <= 'h0;
		'h52 : r_sqroot <= 'h0;
		'h53 : r_sqroot <= 'h0;
		'h54 : r_sqroot <= 'h1;
		'h55 : r_sqroot <= 'h1;
		'h56 : r_sqroot <= 'h1;
		'h57 : r_sqroot <= 'h1;
		'h58 : r_sqroot <= 'h1;
		'h59 : r_sqroot <= 'h2;
		'h5a : r_sqroot <= 'h2;
		'h5b : r_sqroot <= 'h2;
		'h5c : r_sqroot <= 'h2;
		'h5d : r_sqroot <= 'h2;
		'h5e : r_sqroot <= 'h3;
		'h5f : r_sqroot <= 'h3;
		'h60 : r_sqroot <= 'h3;
		'h61 : r_sqroot <= 'h3;
		'h62 : r_sqroot <= 'h3;
		'h63 : r_sqroot <= 'h4;
		'h64 : r_sqroot <= 'h4;
		'h65 : r_sqroot <= 'h4;
		'h66 : r_sqroot <= 'h4;
		'h67 : r_sqroot <= 'h4;
		'h68 : r_sqroot <= 'h4;
		'h69 : r_sqroot <= 'h5;
		'h6a : r_sqroot <= 'h5;
		'h6b : r_sqroot <= 'h5;
		'h6c : r_sqroot <= 'h5;
		'h6d : r_sqroot <= 'h5;
		'h6e : r_sqroot <= 'h5;
		'h6f : r_sqroot <= 'h6;
		'h70 : r_sqroot <= 'h6;
		'h71 : r_sqroot <= 'h6;
		'h72 : r_sqroot <= 'h6;
		'h73 : r_sqroot <= 'h6;
		'h74 : r_sqroot <= 'h6;
		'h75 : r_sqroot <= 'h7;
		'h76 : r_sqroot <= 'h7;
		'h77 : r_sqroot <= 'h7;
		'h78 : r_sqroot <= 'h7;
		'h79 : r_sqroot <= 'h7;
		'h7a : r_sqroot <= 'h7;
		'h7b : r_sqroot <= 'h8;
		'h7c : r_sqroot <= 'h8;
		'h7d : r_sqroot <= 'h8;
		'h7e : r_sqroot <= 'h8;
		'h7f : r_sqroot <= 'h8;
		'h80 : r_sqroot <= 'h8;
		'h81 : r_sqroot <= 'h9;
		'h82 : r_sqroot <= 'h9;
		'h83 : r_sqroot <= 'h9;
		'h84 : r_sqroot <= 'h9;
		'h85 : r_sqroot <= 'h9;
		'h86 : r_sqroot <= 'h9;
		'h87 : r_sqroot <= 'ha;
		'h88 : r_sqroot <= 'ha;
		'h89 : r_sqroot <= 'ha;
		'h8a : r_sqroot <= 'ha;
		'h8b : r_sqroot <= 'ha;
		'h8c : r_sqroot <= 'ha;
		'h8d : r_sqroot <= 'ha;
		'h8e : r_sqroot <= 'hb;
		'h8f : r_sqroot <= 'hb;
		'h90 : r_sqroot <= 'hb;
		'h91 : r_sqroot <= 'hb;
		'h92 : r_sqroot <= 'hb;
		'h93 : r_sqroot <= 'hb;
		'h94 : r_sqroot <= 'hc;
		'h95 : r_sqroot <= 'hc;
		'h96 : r_sqroot <= 'hc;
		'h97 : r_sqroot <= 'hc;
		'h98 : r_sqroot <= 'hc;
		'h99 : r_sqroot <= 'hc;
		'h9a : r_sqroot <= 'hc;
		'h9b : r_sqroot <= 'hd;
		'h9c : r_sqroot <= 'hd;
		'h9d : r_sqroot <= 'hd;
		'h9e : r_sqroot <= 'hd;
		'h9f : r_sqroot <= 'hd;
		'ha0 : r_sqroot <= 'hd;
		'ha1 : r_sqroot <= 'hd;
		'ha2 : r_sqroot <= 'he;
		'ha3 : r_sqroot <= 'he;
		'ha4 : r_sqroot <= 'he;
		'ha5 : r_sqroot <= 'he;
		'ha6 : r_sqroot <= 'he;
		'ha7 : r_sqroot <= 'he;
		'ha8 : r_sqroot <= 'he;
		'ha9 : r_sqroot <= 'hf;
		'haa : r_sqroot <= 'hf;
		'hab : r_sqroot <= 'hf;
		'hac : r_sqroot <= 'hf;
		'had : r_sqroot <= 'hf;
		'hae : r_sqroot <= 'hf;
		'haf : r_sqroot <= 'hf;
		'hb0 : r_sqroot <= 'h0;
		'hb1 : r_sqroot <= 'h0;
		'hb2 : r_sqroot <= 'h0;
		'hb3 : r_sqroot <= 'h0;
		'hb4 : r_sqroot <= 'h0;
		'hb5 : r_sqroot <= 'h0;
		'hb6 : r_sqroot <= 'h0;
		'hb7 : r_sqroot <= 'h0;
		'hb8 : r_sqroot <= 'h1;
		'hb9 : r_sqroot <= 'h1;
		'hba : r_sqroot <= 'h1;
		'hbb : r_sqroot <= 'h1;
		'hbc : r_sqroot <= 'h1;
		'hbd : r_sqroot <= 'h1;
		'hbe : r_sqroot <= 'h1;
		'hbf : r_sqroot <= 'h2;
		'hc0 : r_sqroot <= 'h2;
		'hc1 : r_sqroot <= 'h2;
		'hc2 : r_sqroot <= 'h2;
		'hc3 : r_sqroot <= 'h2;
		'hc4 : r_sqroot <= 'h2;
		'hc5 : r_sqroot <= 'h2;
		'hc6 : r_sqroot <= 'h2;
		'hc7 : r_sqroot <= 'h3;
		'hc8 : r_sqroot <= 'h3;
		'hc9 : r_sqroot <= 'h3;
		'hca : r_sqroot <= 'h3;
		'hcb : r_sqroot <= 'h3;
		'hcc : r_sqroot <= 'h3;
		'hcd : r_sqroot <= 'h3;
		'hce : r_sqroot <= 'h3;
		'hcf : r_sqroot <= 'h4;
		'hd0 : r_sqroot <= 'h4;
		'hd1 : r_sqroot <= 'h4;
		'hd2 : r_sqroot <= 'h4;
		'hd3 : r_sqroot <= 'h4;
		'hd4 : r_sqroot <= 'h4;
		'hd5 : r_sqroot <= 'h4;
		'hd6 : r_sqroot <= 'h4;
		'hd7 : r_sqroot <= 'h5;
		'hd8 : r_sqroot <= 'h5;
		'hd9 : r_sqroot <= 'h5;
		'hda : r_sqroot <= 'h5;
		'hdb : r_sqroot <= 'h5;
		'hdc : r_sqroot <= 'h5;
		'hdd : r_sqroot <= 'h5;
		'hde : r_sqroot <= 'h5;
		'hdf : r_sqroot <= 'h6;
		'he0 : r_sqroot <= 'h6;
		'he1 : r_sqroot <= 'h6;
		'he2 : r_sqroot <= 'h6;
		'he3 : r_sqroot <= 'h6;
		'he4 : r_sqroot <= 'h6;
		'he5 : r_sqroot <= 'h6;
		'he6 : r_sqroot <= 'h6;
		'he7 : r_sqroot <= 'h7;
		'he8 : r_sqroot <= 'h7;
		'he9 : r_sqroot <= 'h7;
		'hea : r_sqroot <= 'h7;
		'heb : r_sqroot <= 'h7;
		'hec : r_sqroot <= 'h7;
		'hed : r_sqroot <= 'h7;
		'hee : r_sqroot <= 'h7;
		'hef : r_sqroot <= 'h7;
		'hf0 : r_sqroot <= 'h8;
		'hf1 : r_sqroot <= 'h8;
		'hf2 : r_sqroot <= 'h8;
		'hf3 : r_sqroot <= 'h8;
		'hf4 : r_sqroot <= 'h8;
		'hf5 : r_sqroot <= 'h8;
		'hf6 : r_sqroot <= 'h8;
		'hf7 : r_sqroot <= 'h8;
		'hf8 : r_sqroot <= 'h9;
		'hf9 : r_sqroot <= 'h9;
		'hfa : r_sqroot <= 'h9;
		'hfb : r_sqroot <= 'h9;
		'hfc : r_sqroot <= 'h9;
		'hfd : r_sqroot <= 'h9;
		'hfe : r_sqroot <= 'h9;
		'hff : r_sqroot <= 'h9;
		'h100 : r_sqroot <= 'h9;
		'h101 : r_sqroot <= 'ha;
		'h102 : r_sqroot <= 'ha;
		'h103 : r_sqroot <= 'ha;
		'h104 : r_sqroot <= 'ha;
		'h105 : r_sqroot <= 'ha;
		'h106 : r_sqroot <= 'ha;
		'h107 : r_sqroot <= 'ha;
		'h108 : r_sqroot <= 'ha;
		'h109 : r_sqroot <= 'ha;
		'h10a : r_sqroot <= 'hb;
		'h10b : r_sqroot <= 'hb;
		'h10c : r_sqroot <= 'hb;
		'h10d : r_sqroot <= 'hb;
		'h10e : r_sqroot <= 'hb;
		'h10f : r_sqroot <= 'hb;
		'h110 : r_sqroot <= 'hb;
		'h111 : r_sqroot <= 'hb;
		'h112 : r_sqroot <= 'hb;
		'h113 : r_sqroot <= 'hc;
		'h114 : r_sqroot <= 'hc;
		'h115 : r_sqroot <= 'hc;
		'h116 : r_sqroot <= 'hc;
		'h117 : r_sqroot <= 'hc;
		'h118 : r_sqroot <= 'hc;
		'h119 : r_sqroot <= 'hc;
		'h11a : r_sqroot <= 'hc;
		'h11b : r_sqroot <= 'hc;
		'h11c : r_sqroot <= 'hd;
		'h11d : r_sqroot <= 'hd;
		'h11e : r_sqroot <= 'hd;
		'h11f : r_sqroot <= 'hd;
		'h120 : r_sqroot <= 'hd;
		'h121 : r_sqroot <= 'hd;
		'h122 : r_sqroot <= 'hd;
		'h123 : r_sqroot <= 'hd;
		'h124 : r_sqroot <= 'hd;
		'h125 : r_sqroot <= 'hd;
		'h126 : r_sqroot <= 'he;
		'h127 : r_sqroot <= 'he;
		'h128 : r_sqroot <= 'he;
		'h129 : r_sqroot <= 'he;
		'h12a : r_sqroot <= 'he;
		'h12b : r_sqroot <= 'he;
		'h12c : r_sqroot <= 'he;
		'h12d : r_sqroot <= 'he;
		'h12e : r_sqroot <= 'he;
		'h12f : r_sqroot <= 'hf;
		'h130 : r_sqroot <= 'hf;
		'h131 : r_sqroot <= 'hf;
		'h132 : r_sqroot <= 'hf;
		'h133 : r_sqroot <= 'hf;
		'h134 : r_sqroot <= 'hf;
		'h135 : r_sqroot <= 'hf;
		'h136 : r_sqroot <= 'hf;
		'h137 : r_sqroot <= 'hf;
		'h138 : r_sqroot <= 'hf;
		default: r_sqroot <= 'h0;
	endcase
end
endmodule
