`default_nettype none
module hypCal (
	input wire [9:0] x_pos,
	input wire [9:0] y_pos,
	input wire clk, rst,
	output reg [4:0] r_sqroot
);
wire [12:0] xy_pos;

wire  [8:0] norm_x = (x_pos[9] == 1'b0) ? x_pos[8:0] : ~(x_pos[8:0]);
wire  [8:0] norm_y = (y_pos[9] == 1'b0) ? y_pos[8:0] : ~(y_pos[8:0]);

reg [6:0]mutlReg;
reg stateCheck;
wire [12:0]multSignal = mutlReg*mutlReg;
reg[12:0] multX, multY;
always @(posedge clk) begin
	if (rst) begin
		mutlReg <= 6'h00;
		stateCheck <= 'b0;
	end else begin
		if (stateCheck == 'b0) begin
			multY <=multSignal;
			mutlReg <= norm_x[8:2];
			stateCheck <= 'b1;
		end else begin
			multX <=multSignal;
			mutlReg <= norm_y[8:2];
			stateCheck <= 'b0;
		end
	end
end
		

//assign xy_pos = (norm_y[8:2]*norm_y[8:2] + norm_x[8:2]*norm_x[8:2]) >> 6;
assign xy_pos = (multX + multY) >> 6;
always @(xy_pos) begin
	case(xy_pos)
		'h00 : r_sqroot <= 'h00;
		'h01 : r_sqroot <= 'h03;
		'h02 : r_sqroot <= 'h05;
		'h03 : r_sqroot <= 'h06;
		'h04 : r_sqroot <= 'h07;
		'h05 : r_sqroot <= 'h08;
		'h06 : r_sqroot <= 'h08;
		'h07 : r_sqroot <= 'h09;
		'h08 : r_sqroot <= 'h0a;
		'h09 : r_sqroot <= 'h0a;
		'h0a : r_sqroot <= 'h0b;
		'h0b : r_sqroot <= 'h0c;
		'h0c : r_sqroot <= 'h0c;
		'h0d : r_sqroot <= 'h0d;
		'h0e : r_sqroot <= 'h0d;
		'h0f : r_sqroot <= 'h0e;
		'h10 : r_sqroot <= 'h0e;
		'h11 : r_sqroot <= 'h0e;
		'h12 : r_sqroot <= 'h0f;
		'h13 : r_sqroot <= 'h0f;
		'h14 : r_sqroot <= 'h10;
		'h15 : r_sqroot <= 'h10;
		'h16 : r_sqroot <= 'h10;
		'h17 : r_sqroot <= 'h11;
		'h18 : r_sqroot <= 'h11;
		'h19 : r_sqroot <= 'h12;
		'h1a : r_sqroot <= 'h12;
		'h1b : r_sqroot <= 'h12;
		'h1c : r_sqroot <= 'h13;
		'h1d : r_sqroot <= 'h13;
		'h1e : r_sqroot <= 'h13;
		'h1f : r_sqroot <= 'h14;
		'h20 : r_sqroot <= 'h14;
		'h21 : r_sqroot <= 'h14;
		'h22 : r_sqroot <= 'h15;
		'h23 : r_sqroot <= 'h15;
		'h24 : r_sqroot <= 'h15;
		'h25 : r_sqroot <= 'h16;
		'h26 : r_sqroot <= 'h16;
		'h27 : r_sqroot <= 'h16;
		'h28 : r_sqroot <= 'h16;
		'h29 : r_sqroot <= 'h17;
		'h2a : r_sqroot <= 'h17;
		'h2b : r_sqroot <= 'h17;
		'h2c : r_sqroot <= 'h18;
		'h2d : r_sqroot <= 'h18;
		'h2e : r_sqroot <= 'h18;
		'h2f : r_sqroot <= 'h18;
		'h30 : r_sqroot <= 'h19;
		'h31 : r_sqroot <= 'h19;
		'h32 : r_sqroot <= 'h19;
		'h33 : r_sqroot <= 'h19;
		'h34 : r_sqroot <= 'h1a;
		'h35 : r_sqroot <= 'h1a;
		'h36 : r_sqroot <= 'h1a;
		'h37 : r_sqroot <= 'h1a;
		'h38 : r_sqroot <= 'h1b;
		'h39 : r_sqroot <= 'h1b;
		'h3a : r_sqroot <= 'h1b;
		'h3b : r_sqroot <= 'h1b;
		'h3c : r_sqroot <= 'h1c;
		'h3d : r_sqroot <= 'h1c;
		'h3e : r_sqroot <= 'h1c;
		'h3f : r_sqroot <= 'h1c;
		'h40 : r_sqroot <= 'h1c;
		'h41 : r_sqroot <= 'h1d;
		'h42 : r_sqroot <= 'h1d;
		'h43 : r_sqroot <= 'h1d;
		'h44 : r_sqroot <= 'h1d;
		'h45 : r_sqroot <= 'h1e;
		'h46 : r_sqroot <= 'h1e;
		'h47 : r_sqroot <= 'h1e;
		'h48 : r_sqroot <= 'h1e;
		'h49 : r_sqroot <= 'h1e;
		'h4a : r_sqroot <= 'h1f;
		'h4b : r_sqroot <= 'h1f;
		'h4c : r_sqroot <= 'h1f;
		'h4d : r_sqroot <= 'h1f;
		'h4e : r_sqroot <= 'h1f;
		'h4f : r_sqroot <= 'h20;
		'h50 : r_sqroot <= 'h20;
		'h51 : r_sqroot <= 'h20;
		'h52 : r_sqroot <= 'h20;
		'h53 : r_sqroot <= 'h20;
		'h54 : r_sqroot <= 'h21;
		'h55 : r_sqroot <= 'h21;
		'h56 : r_sqroot <= 'h21;
		'h57 : r_sqroot <= 'h21;
		'h58 : r_sqroot <= 'h21;
		'h59 : r_sqroot <= 'h22;
		'h5a : r_sqroot <= 'h22;
		'h5b : r_sqroot <= 'h22;
		'h5c : r_sqroot <= 'h22;
		'h5d : r_sqroot <= 'h22;
		'h5e : r_sqroot <= 'h23;
		'h5f : r_sqroot <= 'h23;
		'h60 : r_sqroot <= 'h23;
		'h61 : r_sqroot <= 'h23;
		'h62 : r_sqroot <= 'h23;
		'h63 : r_sqroot <= 'h24;
		'h64 : r_sqroot <= 'h24;
		'h65 : r_sqroot <= 'h24;
		'h66 : r_sqroot <= 'h24;
		'h67 : r_sqroot <= 'h24;
		'h68 : r_sqroot <= 'h24;
		'h69 : r_sqroot <= 'h25;
		'h6a : r_sqroot <= 'h25;
		'h6b : r_sqroot <= 'h25;
		'h6c : r_sqroot <= 'h25;
		'h6d : r_sqroot <= 'h25;
		'h6e : r_sqroot <= 'h25;
		'h6f : r_sqroot <= 'h26;
		'h70 : r_sqroot <= 'h26;
		'h71 : r_sqroot <= 'h26;
		'h72 : r_sqroot <= 'h26;
		'h73 : r_sqroot <= 'h26;
		'h74 : r_sqroot <= 'h26;
		'h75 : r_sqroot <= 'h27;
		'h76 : r_sqroot <= 'h27;
		'h77 : r_sqroot <= 'h27;
		'h78 : r_sqroot <= 'h27;
		'h79 : r_sqroot <= 'h27;
		'h7a : r_sqroot <= 'h27;
		'h7b : r_sqroot <= 'h28;
		'h7c : r_sqroot <= 'h28;
		'h7d : r_sqroot <= 'h28;
		'h7e : r_sqroot <= 'h28;
		'h7f : r_sqroot <= 'h28;
		'h80 : r_sqroot <= 'h28;
		'h81 : r_sqroot <= 'h29;
		'h82 : r_sqroot <= 'h29;
		'h83 : r_sqroot <= 'h29;
		'h84 : r_sqroot <= 'h29;
		'h85 : r_sqroot <= 'h29;
		'h86 : r_sqroot <= 'h29;
		'h87 : r_sqroot <= 'h2a;
		'h88 : r_sqroot <= 'h2a;
		'h89 : r_sqroot <= 'h2a;
		'h8a : r_sqroot <= 'h2a;
		'h8b : r_sqroot <= 'h2a;
		'h8c : r_sqroot <= 'h2a;
		'h8d : r_sqroot <= 'h2a;
		'h8e : r_sqroot <= 'h2b;
		'h8f : r_sqroot <= 'h2b;
		'h90 : r_sqroot <= 'h2b;
		'h91 : r_sqroot <= 'h2b;
		'h92 : r_sqroot <= 'h2b;
		'h93 : r_sqroot <= 'h2b;
		'h94 : r_sqroot <= 'h2c;
		'h95 : r_sqroot <= 'h2c;
		'h96 : r_sqroot <= 'h2c;
		'h97 : r_sqroot <= 'h2c;
		'h98 : r_sqroot <= 'h2c;
		'h99 : r_sqroot <= 'h2c;
		'h9a : r_sqroot <= 'h2c;
		'h9b : r_sqroot <= 'h2d;
		'h9c : r_sqroot <= 'h2d;
		'h9d : r_sqroot <= 'h2d;
		'h9e : r_sqroot <= 'h2d;
		'h9f : r_sqroot <= 'h2d;
		'ha0 : r_sqroot <= 'h2d;
		'ha1 : r_sqroot <= 'h2d;
		'ha2 : r_sqroot <= 'h2e;
		'ha3 : r_sqroot <= 'h2e;
		'ha4 : r_sqroot <= 'h2e;
		'ha5 : r_sqroot <= 'h2e;
		'ha6 : r_sqroot <= 'h2e;
		'ha7 : r_sqroot <= 'h2e;
		'ha8 : r_sqroot <= 'h2e;
		'ha9 : r_sqroot <= 'h2f;
		'haa : r_sqroot <= 'h2f;
		'hab : r_sqroot <= 'h2f;
		'hac : r_sqroot <= 'h2f;
		'had : r_sqroot <= 'h2f;
		'hae : r_sqroot <= 'h2f;
		'haf : r_sqroot <= 'h2f;
		'hb0 : r_sqroot <= 'h30;
		'hb1 : r_sqroot <= 'h30;
		'hb2 : r_sqroot <= 'h30;
		'hb3 : r_sqroot <= 'h30;
		'hb4 : r_sqroot <= 'h30;
		'hb5 : r_sqroot <= 'h30;
		'hb6 : r_sqroot <= 'h30;
		'hb7 : r_sqroot <= 'h30;
		'hb8 : r_sqroot <= 'h31;
		'hb9 : r_sqroot <= 'h31;
		'hba : r_sqroot <= 'h31;
		'hbb : r_sqroot <= 'h31;
		'hbc : r_sqroot <= 'h31;
		'hbd : r_sqroot <= 'h31;
		'hbe : r_sqroot <= 'h31;
		'hbf : r_sqroot <= 'h32;
		'hc0 : r_sqroot <= 'h32;
		'hc1 : r_sqroot <= 'h32;
		'hc2 : r_sqroot <= 'h32;
		'hc3 : r_sqroot <= 'h32;
		'hc4 : r_sqroot <= 'h32;
		'hc5 : r_sqroot <= 'h32;
		'hc6 : r_sqroot <= 'h32;
		'hc7 : r_sqroot <= 'h33;
		'hc8 : r_sqroot <= 'h33;
		'hc9 : r_sqroot <= 'h33;
		'hca : r_sqroot <= 'h33;
		'hcb : r_sqroot <= 'h33;
		'hcc : r_sqroot <= 'h33;
		'hcd : r_sqroot <= 'h33;
		'hce : r_sqroot <= 'h33;
		'hcf : r_sqroot <= 'h34;
		'hd0 : r_sqroot <= 'h34;
		'hd1 : r_sqroot <= 'h34;
		'hd2 : r_sqroot <= 'h34;
		'hd3 : r_sqroot <= 'h34;
		'hd4 : r_sqroot <= 'h34;
		'hd5 : r_sqroot <= 'h34;
		'hd6 : r_sqroot <= 'h34;
		'hd7 : r_sqroot <= 'h35;
		'hd8 : r_sqroot <= 'h35;
		'hd9 : r_sqroot <= 'h35;
		'hda : r_sqroot <= 'h35;
		'hdb : r_sqroot <= 'h35;
		'hdc : r_sqroot <= 'h35;
		'hdd : r_sqroot <= 'h35;
		'hde : r_sqroot <= 'h35;
		'hdf : r_sqroot <= 'h36;
		'he0 : r_sqroot <= 'h36;
		'he1 : r_sqroot <= 'h36;
		'he2 : r_sqroot <= 'h36;
		'he3 : r_sqroot <= 'h36;
		'he4 : r_sqroot <= 'h36;
		'he5 : r_sqroot <= 'h36;
		'he6 : r_sqroot <= 'h36;
		'he7 : r_sqroot <= 'h37;
		'he8 : r_sqroot <= 'h37;
		'he9 : r_sqroot <= 'h37;
		'hea : r_sqroot <= 'h37;
		'heb : r_sqroot <= 'h37;
		'hec : r_sqroot <= 'h37;
		'hed : r_sqroot <= 'h37;
		'hee : r_sqroot <= 'h37;
		'hef : r_sqroot <= 'h37;
		'hf0 : r_sqroot <= 'h38;
		'hf1 : r_sqroot <= 'h38;
		'hf2 : r_sqroot <= 'h38;
		'hf3 : r_sqroot <= 'h38;
		'hf4 : r_sqroot <= 'h38;
		'hf5 : r_sqroot <= 'h38;
		'hf6 : r_sqroot <= 'h38;
		'hf7 : r_sqroot <= 'h38;
		'hf8 : r_sqroot <= 'h39;
		'hf9 : r_sqroot <= 'h39;
		'hfa : r_sqroot <= 'h39;
		'hfb : r_sqroot <= 'h39;
		'hfc : r_sqroot <= 'h39;
		'hfd : r_sqroot <= 'h39;
		'hfe : r_sqroot <= 'h39;
		'hff : r_sqroot <= 'h39;
		'h100 : r_sqroot <= 'h39;
		'h101 : r_sqroot <= 'h3a;
		'h102 : r_sqroot <= 'h3a;
		'h103 : r_sqroot <= 'h3a;
		'h104 : r_sqroot <= 'h3a;
		'h105 : r_sqroot <= 'h3a;
		'h106 : r_sqroot <= 'h3a;
		'h107 : r_sqroot <= 'h3a;
		'h108 : r_sqroot <= 'h3a;
		'h109 : r_sqroot <= 'h3a;
		'h10a : r_sqroot <= 'h3b;
		'h10b : r_sqroot <= 'h3b;
		'h10c : r_sqroot <= 'h3b;
		'h10d : r_sqroot <= 'h3b;
		'h10e : r_sqroot <= 'h3b;
		'h10f : r_sqroot <= 'h3b;
		'h110 : r_sqroot <= 'h3b;
		'h111 : r_sqroot <= 'h3b;
		'h112 : r_sqroot <= 'h3b;
		'h113 : r_sqroot <= 'h3c;
		'h114 : r_sqroot <= 'h3c;
		'h115 : r_sqroot <= 'h3c;
		'h116 : r_sqroot <= 'h3c;
		'h117 : r_sqroot <= 'h3c;
		'h118 : r_sqroot <= 'h3c;
		'h119 : r_sqroot <= 'h3c;
		'h11a : r_sqroot <= 'h3c;
		'h11b : r_sqroot <= 'h3c;
		'h11c : r_sqroot <= 'h3d;
		'h11d : r_sqroot <= 'h3d;
		'h11e : r_sqroot <= 'h3d;
		'h11f : r_sqroot <= 'h3d;
		'h120 : r_sqroot <= 'h3d;
		'h121 : r_sqroot <= 'h3d;
		'h122 : r_sqroot <= 'h3d;
		'h123 : r_sqroot <= 'h3d;
		'h124 : r_sqroot <= 'h3d;
		'h125 : r_sqroot <= 'h3d;
		'h126 : r_sqroot <= 'h3e;
		'h127 : r_sqroot <= 'h3e;
		'h128 : r_sqroot <= 'h3e;
		'h129 : r_sqroot <= 'h3e;
		'h12a : r_sqroot <= 'h3e;
		'h12b : r_sqroot <= 'h3e;
		'h12c : r_sqroot <= 'h3e;
		'h12d : r_sqroot <= 'h3e;
		'h12e : r_sqroot <= 'h3e;
		'h12f : r_sqroot <= 'h3f;
		'h130 : r_sqroot <= 'h3f;
		'h131 : r_sqroot <= 'h3f;
		'h132 : r_sqroot <= 'h3f;
		'h133 : r_sqroot <= 'h3f;
		'h134 : r_sqroot <= 'h3f;
		'h135 : r_sqroot <= 'h3f;
		'h136 : r_sqroot <= 'h3f;
		'h137 : r_sqroot <= 'h3f;
		'h138 : r_sqroot <= 'h3f;
		default: r_sqroot <= 'h00;
	endcase
end
endmodule
